library ieee;
use ieee.std_logic_1164.all;

entity alu is
    port (
      clock    : in    std_logic;       
      reset    : in    std_logic;       
      cpu_bus  : inout std_logic_vector(31 downto 0);  
      s_code   : in    std_logic_vector(11 downto 0);  
      a_in     : in    std_logic;       
      c_in     : in    std_logic;       
      c_out    : in    std_logic       
      );
end alu;

architecture rtl of alu is

component A_register is
  port (
    clock : in  std_logic;              
    reset : in  std_logic;              
    d     : in  std_logic_vector(31 downto 0);  
    q     : out std_logic_vector(31 downto 0);  
    load  : in  std_logic               
    );
end component;


  component C_register is
  port (
    clock   : in  std_logic;           
    reset   : in  std_logic;           
    d       : in  std_logic_vector(31 downto 0);  
    out_bus : out std_logic_vector(31 downto 0);  
    load    : in  std_logic;            
    E      : in  std_logic             
    );
  end component;
  
  component R_shift is
    port (
      B          : in  std_logic_vector(31 downto 0);  
      C          : out std_logic_vector(31 downto 0);  
      ArthM		  : in  std_logic;       
      Rshift     : in  std_logic        
      );
   end component;

  component L_shift is
    port (
      B          : in  std_logic_vector(31 downto 0);  
      C          : out std_logic_vector(31 downto 0);  
      Cr		     : in  std_logic;       
      Lshift     : in  std_logic        
      );
  end component;

  component adderALU is
  port (
    a    : in  std_logic_vector(31 downto 0);  
    b    : in  std_logic_vector(31 downto 0);  
    c    : out std_logic_vector(31 downto 0); 
    inc4 : in  std_logic;             
    add  : in  std_logic;               
    sub  : in  std_logic;               
    pass : in  std_logic;               
    inv  : in  std_logic;
    neg  : in  std_logic	 
    );
  end component;


 component logic_gate is
  port (
    a           : in  std_logic_vector(31 downto 0);  
    b           : in  std_logic_vector(31 downto 0);  
    c           : out std_logic_vector(31 downto 0);  
    OP_or  		 : in  std_logic;       
    OP_and		 : in  std_logic         
    );
 end component;

  signal s_add    : std_logic ;
  signal s_and    : std_logic ;
  signal s_c_eq_b : std_logic ;
  signal s_inc_4  : std_logic ;
  signal s_not    : std_logic ;
  signal s_or     : std_logic ;
  signal s_sub    : std_logic ;
  signal s_shc    : std_logic ;
  signal s_shl    : std_logic ;
  signal s_shr    : std_logic ;
  signal s_shra   : std_logic ;
  signal s_neg   : std_logic ;

  signal a : std_logic_vector(31 downto 0);

  signal c : std_logic_vector(31 downto 0);
  
begin  


 s_add    <= s_code(0);
 s_and    <= s_code(1); 
 s_c_eq_b <= s_code(2);
 s_inc_4  <= s_code(3);
 s_not    <= s_code(4);
 s_or     <= s_code(5);
 s_sub    <= s_code(6);
 s_shc    <= s_code(7);
 s_shl    <= s_code(8);
 s_shr    <= s_code(9);
 s_shra   <= s_code(10);
 s_neg    <= s_code(11);

  regA      : A_register port map ( clock, reset, cpu_bus, a, a_in );
  regC      : C_register port map ( clock, reset, c , cpu_bus, c_in, c_out );
  r_s       : R_shift    port map ( cpu_bus, c, s_shra, s_shr );
  l_s       : L_shift    port map ( cpu_bus, c, s_shc, s_shl );
  add       : adderALU   port map ( a, cpu_bus, c, s_inc_4, s_add,
                                      s_sub, s_c_eq_b, s_not,s_neg  );
  a_b_AndOR : logic_gate  port map ( a, cpu_bus, c, s_or, s_and );

end rtl;