library ieee;
use ieee.std_logic_1164.all;

entity CPU is
  port (
    master_clock : in    std_logic;     
    start        : in    std_logic;     
    reset        : in    std_logic;    
    done         : in    std_logic;    
    md_read      : in    std_logic;   
    md_write     : in    std_logic;    
    r            : out   std_logic;    
    w            : out   std_logic;     
    ma           : out   std_logic_vector(31 downto 0);
    md           : inout std_logic_vector(31 downto 0)   
  );
end CPU;



architecture rtl of CPU is

  component control_unit is
  port (
			Master_clock : in std_logic;
		reset			 : in std_logic;
		start 		 : in std_logic;
		
		done  		 : in std_logic;
		
		con   : in std_logic;
		Nzero : in std_logic;
		
		opcode: in std_logic_vector(4 downto 0);

		CONin : OUT std_logic;          
		Rin   : OUT std_logic;
		Rout  : OUT std_logic;
		BAout : OUT std_logic;
		Gra   : OUT std_logic;
		Grb   : OUT std_logic;
		Grc   : OUT std_logic;
		Dec   : OUT std_logic;
		load  : OUT std_logic;          
		C1out : OUT std_logic;
		C2out : OUT std_logic;          
		PCin  : OUT std_logic;
		PCout : OUT std_logic;
		Ain   : OUT std_logic;
		IRin  : OUT std_logic;
		MDin  : OUT std_logic;
		MDout : OUT std_logic;
		MAin  : OUT std_logic;
		Cout  : OUT std_logic;
		Cin   : OUT std_logic;
		
		r     : out std_logic;
		w     : out std_logic;
		
		Add   : OUT std_logic;
		andOp : OUT std_logic;
		CB    : OUT std_logic;
		INC4  : OUT std_logic;
		NOTOP : OUT std_logic;
		OrOP  : OUT std_logic;
		Sub   : OUT std_logic;
		SHC   : OUT std_logic;
		SHL   : OUT std_logic;
		SHR   : OUT std_logic;
		SHRA  : OUT std_logic;
		NEG   : OUT std_logic
		
  );
end component;

component data_path is
  port (
    clock       : in    std_logic;     
    reset       : in    std_logic;     
    r_out       : in    std_logic;      
    r_in        : in    std_logic;    
    g_ra        : in    std_logic;    
    g_rb        : in    std_logic;     
    g_rc        : in    std_logic;      
    ba_out      : in    std_logic;     
    a_in        : in    std_logic;      
    c_in        : in    std_logic;     
    c_out       : in    std_logic;     
    alu_code    : in    std_logic_vector(11 downto 0); 
    pc_out      : in    std_logic;     
    pc_in       : in    std_logic;      
    con         : out   std_logic;     
    con_in      : in    std_logic;     
    c1_out      : in    std_logic;      
    c2_out      : in    std_logic;      
    ir_in       : in    std_logic;     
    opcode      : out   std_logic_vector(4 downto 0); 
    ma          : out   std_logic_vector(31 downto 0);  
    md          : inout std_logic_vector(31 downto 0);  
    ma_in       : in    std_logic;      
    md_bus      : in    std_logic;      
    md_read     : in    std_logic;    
    md_write    : in    std_logic;      
    md_out      : in    std_logic;     
    n_equ_zero  : out   std_logic;     
    n_decrement : in    std_logic;     
    load        : in    std_logic       
    );
end component;

  signal r_out       : std_logic;
 
  signal r_in        : std_logic;
  signal g_ra        : std_logic;
  signal g_rb        : std_logic;
  signal g_rc        : std_logic;
  signal ba_out      : std_logic;
  signal a_in        : std_logic;
  signal c_in        : std_logic;
  signal c_out       : std_logic;
  signal alu_code    : std_logic_vector(11 downto 0);
  signal pc_out      : std_logic;
  signal pc_in       : std_logic;
  signal con         : std_logic;
  signal con_in      : std_logic;
  signal c1_out      : std_logic;
  signal c2_out      : std_logic;
  signal ir_in       : std_logic;
  signal opcode      : std_logic_vector(4 downto 0);
  signal ma_in       : std_logic;
  signal md_in       : std_logic;
  signal md_out      : std_logic;
  signal n_equ_zero  : std_logic;
  signal n_decrement : std_logic;
  signal load        : std_logic;
begin  

  cu : control_unit port map ( master_clock, reset , start, done, con, n_equ_zero,
                               opcode, con_in, r_in, r_out, ba_out, g_ra, g_rb,
                               g_rc , n_decrement, load, c1_out, c2_out, pc_in,
                               pc_out, a_in, ir_in, md_in, md_out, ma_in,
                               c_out, c_in, r, w, alu_code(0),alu_code(1),
										 alu_code(2),alu_code(3),alu_code(4),alu_code(5),
										 alu_code(6),alu_code(7),alu_code(8),alu_code(9),
										 alu_code(10),alu_code(11));
										 
  dp : data_path port map ( master_clock, reset, r_out, r_in, g_ra, g_rb, g_rc,
                            ba_out, a_in, c_in, c_out, alu_code, pc_out, pc_in,
                            con, con_in, c1_out, c2_out, ir_in, opcode, ma,
                            md, ma_in, md_in, md_read, md_write, md_out,
                            n_equ_zero, n_decrement,load );

end rtl;
