library ieee;
use ieee.std_logic_1164.all;

entity shift_counter is
  port (
    clock       : in  std_logic;       
    reset       : in  std_logic;       
    cpu_bus     : in  std_logic_vector(4 downto 0);  
    n_decrement : in  std_logic;       
    n_in        : in  std_logic;       
    n_equ_zero  : out std_logic        
    );
end shift_counter;

architecture rtl of shift_counter is
 
  component D_Flip_Flop
    port (
      clock : in  std_logic;
      reset : in  std_logic;
      d     : in  std_logic;
      q     : out std_logic
      );
  end component;

  signal n   : std_logic_vector(4 downto 0);
  signal sop : std_logic_vector(4 downto 0);
  signal mux : std_logic_vector(4 downto 0);
  
begin  

  sop(0) <=   not n(0);
  
  sop(1) <= ((not n(0)) and (not n(1))) or  (n(0) and n(1));
  
  sop(2) <= ((not n(0)) and (not n(1))  and (not n(2))) or (n(0) and n(2)) 
				or (n(1) and n(2));
				
  sop(3) <= ((not n(0)) and (not n(1)) and (not n(2)) and (not n(3)))
				or (n(0) and n(3))  or (n(1) and n(3)) or (n(2) and n(3));
				
  sop(4) <= ((not n(0)) and (not n(1)) and (not n(2)) and (not n(3)) 
				 and (not n(4)))or (n(0) and n(4)) or (n(1) and n(4))
				or (n(2) and n(4)) or (n(3) and n(4));

process (cpu_bus, sop, n_in, n_decrement,n)
  begin  
    for i in 0 to 4 loop
      mux(i) <= (cpu_bus(i) and n_in)
        or (sop(i) and (not n_in) and n_decrement)
        or (n(i) and (not n_in) and (not n_decrement));
    end loop;  
end process;
  
  dff0 : D_Flip_Flop port map ( clock, reset, mux(0), n(0) );
  dff1 : D_Flip_Flop port map ( clock, reset, mux(1), n(1) );
  dff2 : D_Flip_Flop port map ( clock, reset, mux(2), n(2) );
  dff3 : D_Flip_Flop port map ( clock, reset, mux(3), n(3) );
  dff4 : D_Flip_Flop port map ( clock, reset, mux(4), n(4) );

  n_equ_zero <= not(n(0) or n(1) or n(2) or n(3) or n(4));
  
end rtl;
