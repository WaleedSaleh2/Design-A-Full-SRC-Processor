library ieee;
use ieee.std_logic_1164.all;

entity data_path is
  port (
    clock       : in    std_logic;     
    reset       : in    std_logic;     
    r_out       : in    std_logic;      
    r_in        : in    std_logic;    
    g_ra        : in    std_logic;    
    g_rb        : in    std_logic;     
    g_rc        : in    std_logic;      
    ba_out      : in    std_logic;     
    a_in        : in    std_logic;      
    c_in        : in    std_logic;     
    c_out       : in    std_logic;     
    alu_code    : in    std_logic_vector(11 downto 0); 
    pc_out      : in    std_logic;     
    pc_in       : in    std_logic;      
    con         : out   std_logic;     
    con_in      : in    std_logic;     
    c1_out      : in    std_logic;      
    c2_out      : in    std_logic;      
    ir_in       : in    std_logic;     
    opcode      : out   std_logic_vector(4 downto 0); 
    ma          : out   std_logic_vector(31 downto 0);  
    md          : inout std_logic_vector(31 downto 0);  
    ma_in       : in    std_logic;      
    md_bus      : in    std_logic;      
    md_read     : in    std_logic;    
    md_write    : in    std_logic;      
    md_out      : in    std_logic;     
    n_equ_zero  : out   std_logic;     
    n_decrement : in    std_logic;     
    load        : in    std_logic
    );
end data_path;


architecture data_path_arch of data_path is

  component register_file
    port (
      clock   : in    std_logic;
      reset   : in    std_logic;
      cpu_bus : inout std_logic_vector(31 downto 0);
      ra      : in    std_logic_vector(4 downto 0);
      rb      : in    std_logic_vector(4 downto 0);
      rc      : in    std_logic_vector(4 downto 0);
      g_ra    : in    std_logic;
      g_rb    : in    std_logic;
      g_rc    : in    std_logic;
      r_in    : in    std_logic;
      r_out   : in    std_logic;
      ba_out  : in    std_logic
      );
  end component;

  component alu
    port (
      clock    : in    std_logic;
      reset    : in    std_logic;
      cpu_bus  : inout std_logic_vector(31 downto 0);
      s_code   : in    std_logic_vector(11 downto 0);
      a_in     : in    std_logic;
      c_in     : in    std_logic;
      c_out    : in    std_logic
      );
  end component;

  component PC
    port (
      clock : in    std_logic;
      reset : in    std_logic;
      d_bus : inout std_logic_vector(31 downto 0);  -- cpu_bus
      PCin  : in    std_logic;                      -- pc_in
      PCout : in    std_logic                       -- pc_out
      );
  end component;

  component condition
    port (
      clock   : in    std_logic;
      reset   : in    std_logic;
      cpu_bus : in std_logic_vector(31 downto 0);
      c3      : in    std_logic_vector(2 downto 0);
      con_in  : in    std_logic;
      con     : out   std_logic
      );
  end component;

  component instruction_register
    port (
      clock   : in    std_logic;
      reset   : in    std_logic;
      cpu_bus : inout std_logic_vector(31 downto 0);
      c1_out  : in    std_logic;
      c2_out  : in    std_logic;
      ir_in   : in    std_logic;
      opcode  : out   std_logic_vector(4 downto 0);
      c3      : inout std_logic_vector(2 downto 0);
      ra      : inout std_logic_vector(4 downto 0);
      rb      : inout std_logic_vector(4 downto 0);
      rc      : inout std_logic_vector(4 downto 0)
      );
  end component;

  component memory_interface
    port (
      clock    : in    std_logic;
      reset    : in    std_logic;
      cpu_bus  : inout std_logic_vector(31 downto 0);
      ma       : out   std_logic_vector(31 downto 0);
      md       : inout std_logic_vector(31 downto 0);
      ma_in    : in    std_logic;
      md_bus   : in    std_logic;
      md_read  : in    std_logic;
      md_write : in    std_logic;
      md_out   : in    std_logic
    );
  end component;

  component shift_counter
    port (
      clock       : in    std_logic;
      reset       : in    std_logic;
      cpu_bus     : in    std_logic_vector(4 downto 0);
      n_decrement : in    std_logic;
      n_in        : in    std_logic;
      n_equ_zero  : out   std_logic
      );
  end component;

  signal cpu_bus : std_logic_vector(31 downto 0);
  signal c3      : std_logic_vector(2 downto 0);
  signal ra      : std_logic_vector(4 downto 0);
  signal rb      : std_logic_vector(4 downto 0);
  signal rc      : std_logic_vector(4 downto 0);
  
  signal pc_Input: std_logic_vector(31 downto 0);
  
begin  

  pc_Input    <= cpu_bus or "00000000000000000000000000000000";
 	
  RegFIleL : register_file        port map (clock,reset,cpu_bus,ra,rb,rc,g_ra,g_rb,g_rc,r_in,r_out,ba_out);
  
  ALUL 	  : alu                  port map (clock,reset,cpu_bus,alu_code,a_in, c_in, c_out);
  
  PCL      : PC					    port map (clock,reset,pc_Input,pc_in,pc_out);
  
  CONDL    : condition            port map (clock,reset,cpu_bus,c3,con_in,con);
  
  IRL      : instruction_register port map (clock,reset,cpu_bus,c1_out,c2_out,ir_in,opcode,c3,ra,rb,rc);
  
  MEML     : memory_interface     port map (clock,reset,cpu_bus,ma, md,ma_in,md_bus,md_read,md_write,md_out);
  
  shLable  : shift_counter        port map (clock,reset,cpu_bus(4 downto 0),n_decrement,load,n_equ_zero);
  
end data_path_arch; 
