library ieee;
use ieee.STD_LOGIC_1164.ALL;

entity Controlunitlogic is
    Port ( 		
   		      T0			: in std_logic;
   		      T1			: in std_logic;
   		      T2			: in std_logic;
					T3			: in std_logic;
					T4			: in std_logic;
					T5			: in std_logic;
					T6			: in std_logic;
					T7			: in std_logic;
					
					Nzero    : in std_logic;
					CON 		: in std_logic;

					AddInst 	: in std_logic;
					AddiInst : in std_logic;
					SubInst 	: in std_logic;
					AndInst 	: in std_logic;
					AndiInst : in std_logic;
					OrInst 	: in std_logic;
					OriInst  : in std_logic;
					notInst	: in std_logic;
					negInst  : in std_logic;
					
					SHRInst 	: in std_logic;
					SHRAInst : in std_logic;
					SHLInst  : in std_logic;
					SHCInst  : in std_logic;
					
					BrInst	: in std_logic;
					BrlInst	: in std_logic;
					
					ldInst	: in std_logic;
					ldrInst	: in std_logic;
					stInst	: in std_logic;
					strInst	: in std_logic;
					laInst	: in std_logic;
					larInst	: in std_logic;
					
					stopInst : in std_logic;
 			 
			      Add   : OUT std_logic;
					Sub   : OUT std_logic;
					andOp : OUT std_logic;
					OrOP  : OUT std_logic;
					SHR   : OUT std_logic;
					SHRA  : OUT std_logic;
					SHL   : OUT std_logic;
					SHC   : OUT std_logic;
					NOTOP : OUT std_logic;
					NEG   : OUT std_logic;
					
					CB    : OUT std_logic;
					INC4  : OUT std_logic;
					CONin : OUT std_logic;          
					Rin   : OUT std_logic;
					Rout  : OUT std_logic;
					BAout : OUT std_logic;
					Gra   : OUT std_logic;
					Grb   : OUT std_logic;
					Grc   : OUT std_logic;
					Dec   : OUT std_logic;
					load  : OUT std_logic;          
					C1out : OUT std_logic;
					C2out : OUT std_logic;          
					PCin  : OUT std_logic;
					PCout : OUT std_logic;
					Ain   : OUT std_logic;
					IRin  : OUT std_logic;
					MDin  : OUT std_logic;
					MDout : OUT std_logic;
					MAin  : OUT std_logic;
					Cout  : OUT std_logic;
					EndSignal : OUT std_logic;
					waitSignal: OUT std_logic;
					Cin   : OUT std_logic;
					ReadD : OUT std_logic;
					WriteD: OUT Std_logic;
					Goto6 : out Std_logic;
					stop  : OUT std_logic
					);
end Controlunitlogic ;

architecture rtl of Controlunitlogic is


begin

Add 	<=(T4 and (AddInst OR AddiInst OR ldInst OR ldrInst OR strInst OR stInst OR laInst OR larInst));
Sub 	<=(T4 and  SubInst);
AndOP <=(T4 and (AndInst OR AndiInst));
Orop 	<=(T4 and (OrInst Or OriInst));
SHR 	<=(T6 and (not Nzero) and SHRInst);
SHRA 	<=(T6 and (not Nzero) and SHRAInst);
SHL 	<=(T6 and (not Nzero) and SHLInst);
SHC 	<=(T6 and (not Nzero) and SHCInst);
NOTOP <=(T3 and  Notinst);
Neg	<=(T3 and  NegInst);
CB 	<=(T5 and (SHRInst OR SHRAInst OR SHLInst OR SHCInst));
INC4 	<=(T0);

CONin <=(T3 and  brInst ) OR 
		  (T4 and  brlInst);

Rin   <=(T5 and (Addinst OR AddiInst Or AndInst OR AndiInst Or OrInst Or oriInst Or subInst OR larInst OR laInst)) OR 
		  (T4 and (NotInst OR NegInst)) OR 
		  (T7 and (ldrInst OR ldInst OR SHRInst OR SHRAInst OR SHLInst OR SHCInst)) OR 
		  (T3 and  BrlInst);  

Rout  <=(T3 and (AddInst Or ANdInst OR SubInst Or ORinst Or AddiInst Or ANdiInst Or ORiinst Or Notinst Or NegInst OR brinst)) Or 
		  (T4 and (AddInst Or ANdInst OR SubInst Or ORinst OR brlInst OR brInst OR (nzero and(SHRInst OR SHRAInst OR SHLInst OR SHCInst ) ))) OR 
		  (T5 and (BrlInst or SHRInst OR SHRAInst OR SHLInst OR SHCInst )) OR
		  (T6 and (strInst OR stInst ));

BAout <=(T3 and (ldInst OR stInst OR laInst));	

Gra   <=(T5 and (Addinst OR AddiInst Or AndInst OR AndiInst Or OrInst Or oriInst Or subInst oR larInst OR laInst)) OR 
		  (T4 and (NotInst Or NegInst)) OR
		  (T3 and (brlInst)) Or
		  (T6 and (strInst OR stInst)) OR
		  (T7 and (ldrInst OR ldInst OR SHRInst OR SHRAInst OR SHLInst OR SHCInst));
		  
Grb   <=(T3 and (Addinst OR AddiInst Or AndInst OR AndiInst Or OrInst Or oriInst Or subInst Or ldinst OR stInst Or laInst)) OR  		  
		  (T4 and (brInst)) OR 
		  (T5 and (brlInst or SHRInst OR SHRAInst OR SHLInst OR SHCInst));
		  
Grc 	<=(T4 and (Addinst Or AndInst Or OrInst Or subInst OR brlInst OR (nzero and(SHRInst OR SHRAInst OR SHLInst OR SHCInst )))) Or 
		  (T3 and (NotInst Or NEgInst OR brInst)) ;

Dec 	<=(T6 and (not nzero and (SHRInst OR SHRAInst OR SHLInst OR SHCInst )));
Goto6 <=(T6 and (not nzero and (SHRInst OR SHRAInst OR SHLInst OR SHCInst ))); 

load  <=(T3 and (SHRInst OR SHRAInst OR SHLInst OR SHCInst )) OR
		  (T4 and (nzero and (SHRInst OR SHRAInst OR SHLInst OR SHCInst )));
 
C1out <=(T4 and (strInst OR ldrInst OR larInst)) OR
		  (T3 and (SHRInst OR SHRAInst OR SHLInst OR SHCInst ));
C2out <=(T4 and (addiInst OR andiInst Or OriInst OR ldInst Or stInst Or laInst));

PCin  <=(T1) OR
		  (T4 and brInst and CON) OR
		  (T5 and BrlInst and CON);
		  
PCout	<=(T0) OR
		  (T3 and (ldrInst Or strInst OR larInst OR brlInst));
		  
Ain   <=(T3 and (AddInst Or ANdInst OR SubInst Or ORinst Or AddiInst Or ANdiInst Or ORiinst OR ldinst OR stinst Or ldrinst OR strInst OR laInst OR larInst));

IRin	<=(T2);

MDin 	<=(T6 and (stInst or StrInst));
MDout <=(T2) Or
		  (T7 and (ldrInst Or ldInst));

ReadD  <=(T1) OR
		   (T6 and (ldInst OR ldrInst));
WriteD <=(T7 and (strInst Or stInst));		

Cin 	 <=(T0) OR
		   (T4 and (AddInst Or ANdInst OR SubInst Or ORinst Or AddiInst Or ANdiInst Or ORiinst Or ldInst OR ldrInst Or laInst Or larInst OR stInst Or StrInst)) OR
			(T3 and (NotInst OR NegInst)) OR
			(T5 and (SHRInst OR SHRAInst OR SHLInst OR SHCInst)) OR
			(T6 and (not nzero and (SHRInst OR SHRAInst OR SHLInst OR SHCInst )));
			
Cout 	 <=(T1) OR
			(T5 and (AddInst Or ANdInst OR SubInst Or ORinst Or AddiInst Or ANdiInst Or ORiinst Or ldInst OR ldrInst Or laInst Or larInst OR stInst Or StrInst)) OR
			(T4 and (NotInst OR NegInst)) OR
			(T6 and (not nzero and (SHRInst OR SHRAInst OR SHLInst OR SHCInst ))) OR
			(T6 and Nzero) ;
			
MAin 	 <=(T0) OR
			(T5 and (ldInst OR StInst Or ldrInst Or StrInst));
			
waitSignal <= T1                      
              or (T6 and ldInst)     
              or (T6 and ldrInst)   
              or (T7 and stInst)     
              or (T7 and strInst);  
				  
stop 		<=  T3 and stopInst;  
 
EndSignal <= (T4 and (NotInst Or NegInst OR brInst)) OR
				 (T5 and (AddInst Or ANdInst OR SubInst Or ORinst Or AddiInst Or ANdiInst Or ORiinst Or brlInst Or laInst OR larInst)) OR
				 (T7 and (stInst Or strInst Or ldInst Or ldrInst Or SHRInst OR SHRAInst OR SHLInst OR SHCInst ));

end rtl;