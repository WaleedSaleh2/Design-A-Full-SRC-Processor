library ieee;
use ieee.std_logic_1164.all;

entity L_shift is
    port (
      B          : in  std_logic_vector(31 downto 0);  
      C          : out std_logic_vector(31 downto 0);  
      Cr 		  : in  std_logic;       
      Lshift     : in  std_logic        
      );
end L_shift;

architecture rtl of L_shift is

component Buffer_32 is
  port (
    input  : in  std_logic_vector(31 downto 0);  
    output : out std_logic_vector(31 downto 0);  
    enable : in  std_logic              
    );
end component;

  signal Eout : std_logic;
  signal shift : std_logic_vector(31 downto 0);
begin 

  Eout <= Cr or Lshift;

  shift <= B(30 downto 0) & (Cr and B(31));

  shift_buff : Buffer_32 port map ( shift, C, Eout );

end rtl;
