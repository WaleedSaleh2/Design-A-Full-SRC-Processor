library ieee;
use ieee.std_logic_1164.all;

entity D_Flip_Flop is
  port (
    clock : in  std_logic;              
    reset : in  std_logic;              
    d     : in  std_logic;              
    q     : out std_logic               
    );
end D_Flip_Flop;

architecture rtl of D_Flip_Flop is

begin  

process (clock, reset, d)
begin  
   if reset = '1' then
     q <= '0';
   elsif rising_edge( clock ) then
     q <= d;
   end if;
end process;

end rtl;
