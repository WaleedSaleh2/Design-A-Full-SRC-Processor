library ieee;
use ieee.std_logic_1164.all;

entity control_unit is
  port (
		Master_clock : in std_logic;
		reset			 : in std_logic;
		start 		 : in std_logic;
		
		done  		 : in std_logic;
		
		con   : in std_logic;
		Nzero : in std_logic;
		
		opcode: in std_logic_vector(4 downto 0);

		CONin : OUT std_logic;          
		Rin   : OUT std_logic;
		Rout  : OUT std_logic;
		BAout : OUT std_logic;
		Gra   : OUT std_logic;
		Grb   : OUT std_logic;
		Grc   : OUT std_logic;
		Dec   : OUT std_logic;
		load  : OUT std_logic;          
		C1out : OUT std_logic;
		C2out : OUT std_logic;          
		PCin  : OUT std_logic;
		PCout : OUT std_logic;
		Ain   : OUT std_logic;
		IRin  : OUT std_logic;
		MDin  : OUT std_logic;
		MDout : OUT std_logic;
		MAin  : OUT std_logic;
		Cout  : OUT std_logic;
		Cin   : OUT std_logic;
		
		r     : out std_logic;
		w     : out std_logic;
		
		Add   : OUT std_logic;
		andOp : OUT std_logic;
		CB    : OUT std_logic;
		INC4  : OUT std_logic;
		NOTOP : OUT std_logic;
		OrOP  : OUT std_logic;
		Sub   : OUT std_logic;
		SHC   : OUT std_logic;
		SHL   : OUT std_logic;
		SHR   : OUT std_logic;
		SHRA  : OUT std_logic;
		NEG   : OUT std_logic
		
  );
end control_unit;

architecture control_unit_arch of control_unit is

component clocking_logic is
  port (
    clock    : in  std_logic;           
    start    : in  std_logic;          
    reset    : in  std_logic;          
    stop     : in  std_logic;           
    cpu_wait : in  std_logic;          
    done     : in  std_logic;          
    enable   : out std_logic;        
    read_m   : in  std_logic;           
    write_m  : in  std_logic;         
    r        : out std_logic;         
    w        : out std_logic           
    );
end component;

component step_generator is
  port (
    clock    : in  std_logic;           
    enable   : in  std_logic;           
    end_inst : in  std_logic;           
    goto6    : in  std_logic;           
    T0out 	 : out std_logic;
	 T1out 	 : out std_logic;
	 T2out 	 : out std_logic;
	 T3out 	 : out std_logic;
	 T4out    : out std_logic;
	 T5out 	 : out std_logic;
	 T6out 	 : out std_logic;
	 T7out 	 : out std_logic
    );
end component;

component op_code_decoder is
  port (
   input    : in  std_logic_vector(4 downto 0);  
   AddInst 	: out std_logic;
	AddiInst : out std_logic;
	SubInst 	: out std_logic;
	AndInst 	: out std_logic;
	AndiInst : out std_logic;
	OrInst 	: out std_logic;
	OriInst  : out std_logic;
	notInst	: out std_logic;
	negInst  : out std_logic;
	SHRInst 	: out std_logic;
	SHRAInst : out std_logic;
	SHLInst  : out std_logic;
	SHCInst  : out std_logic;
	BrInst	: out std_logic;
	BrlInst	: out std_logic;
	ldInst	: out std_logic;
	ldrInst	: out std_logic;
	stInst	: out std_logic;
	strInst	: out std_logic;
	laInst	: out std_logic;
	larInst	: out std_logic;
	stopInst : out std_logic

	);
end component;

component Controlunitlogic is
    Port ( 		
   		      T0			: in std_logic;
   		      T1			: in std_logic;
   		      T2			: in std_logic;
					T3			: in std_logic;
					T4			: in std_logic;
					T5			: in std_logic;
					T6			: in std_logic;
					T7			: in std_logic;
					
					Nzero    : in std_logic;
					CON 		: in std_logic;

					AddInst 	: in std_logic;
					AddiInst : in std_logic;
					SubInst 	: in std_logic;
					AndInst 	: in std_logic;
					AndiInst : in std_logic;
					OrInst 	: in std_logic;
					OriInst  : in std_logic;
					notInst	: in std_logic;
					negInst  : in std_logic;
					
					SHRInst 	: in std_logic;
					SHRAInst : in std_logic;
					SHLInst  : in std_logic;
					SHCInst  : in std_logic;
					
					BrInst	: in std_logic;
					BrlInst	: in std_logic;
					
					ldInst	: in std_logic;
					ldrInst	: in std_logic;
					stInst	: in std_logic;
					strInst	: in std_logic;
					laInst	: in std_logic;
					larInst	: in std_logic;
					
					stopInst : in std_logic;
 			 
			      Add   : OUT std_logic;
					Sub   : OUT std_logic;
					andOp : OUT std_logic;
					OrOP  : OUT std_logic;
					SHR   : OUT std_logic;
					SHRA  : OUT std_logic;
					SHL   : OUT std_logic;
					SHC   : OUT std_logic;
					NOTOP : OUT std_logic;
					NEG   : OUT std_logic;
					
					CB    : OUT std_logic;
					INC4  : OUT std_logic;
					CONin : OUT std_logic;          
					Rin   : OUT std_logic;
					Rout  : OUT std_logic;
					BAout : OUT std_logic;
					Gra   : OUT std_logic;
					Grb   : OUT std_logic;
					Grc   : OUT std_logic;
					Dec   : OUT std_logic;
					load  : OUT std_logic;          
					C1out : OUT std_logic;
					C2out : OUT std_logic;          
					PCin  : OUT std_logic;
					PCout : OUT std_logic;
					Ain   : OUT std_logic;
					IRin  : OUT std_logic;
					MDin  : OUT std_logic;
					MDout : OUT std_logic;
					MAin  : OUT std_logic;
					Cout  : OUT std_logic;
					EndSignal : OUT std_logic;
					waitSignal: OUT std_logic;
					Cin   : OUT std_logic;
					ReadD : OUT std_logic;
					WriteD: OUT Std_logic;
					Goto6 : out Std_logic;
					stop  : out std_logic
					);
end component;
   
  signal enable    :  std_logic;
  signal sigT0out,
			sigT1out,
			sigT2out,
			sigT3out,
			sigT4out,
			sigT5out,
			sigT6out,
			sigT7out  :  std_logic;
  
   signal cpu_wait :  std_logic;
   signal stop     :  std_logic;
   signal goto6    :  std_logic;
   signal end_inst :  std_logic;
   signal read_m   :  std_logic;
   signal write_m  :  std_logic;
  
   signal AddInst  :  std_logic;
   signal AddiInst :  std_logic;
   signal SubInst  :  std_logic;
	signal AndInst  :  std_logic;
	signal AndiInst :  std_logic;
	signal OrInst 	 :  std_logic;
	signal OriInst  :  std_logic;
	signal notInst	 :  std_logic;
	signal negInst  :  std_logic;
	signal SHRInst  :  std_logic;
	signal SHRAInst :  std_logic;
	signal SHLInst  :  std_logic;
	signal SHCInst  :  std_logic;
	signal BrInst	 :  std_logic;
	signal BrlInst	 :  std_logic;
	signal ldInst	 :  std_logic;
	signal ldrInst	 :  std_logic;
	signal stInst	 :  std_logic;
	signal strInst	 :  std_logic;
	signal laInst	 :  std_logic;
	signal larInst	 :  std_logic;
	signal stopInst :  std_logic;
  
begin  
	 
st: step_generator port map (
  Master_clock,
  enable 	  ,
  end_inst	  ,
  goto6 		  ,
  sigT0out	  ,
  sigT1out 	  ,
  sigT2out 	  ,
  sigT3out 	  ,
  sigT4out 	  ,
  sigT5out 	  ,
  sigT6out 	  ,
  sigT7out 	  
);
  
clock_logic: clocking_logic port map (
  Master_clock ,
  start 			,
  reset 			,
  stop 			, 
  cpu_wait 		,
  done 			, 
  enable 		, 
  read_m 		, 
  write_m 		,
  r 				, 
  w 				
);

de: op_code_decoder port map (
  opcode 		,
  AddInst 		,  
  AddiInst 		, 
  SubInst 		,
  AndInst 		, 
  AndiInst 		, 
  OrInst 		,   
  OriInst 		,
  notInst 		, 
  negInst 		,  
  SHRInst 		,  
  SHRAInst 		,
  SHLInst 		, 
  SHCInst 		, 
  BrInst 		,  
  BrlInst 		, 
  ldInst 		, 
  ldrInst 		, 
  stInst 		,  
  strInst 		,
  laInst 		, 
  larInst 		,
  stopInst
);
	
control: Controlunitlogic port map 
(
sigT0out  ,
sigT1out  ,
sigT2out  ,
sigT3out  ,
sigT4out  ,
sigT5out  ,
sigT6out  ,
sigT7out  ,
Nzero     ,
con       ,
AddInst   ,
AddiInst  ,
SubInst   ,
AndInst   , 
AndiInst  , 
OrInst    ,   
OriInst   ,
notInst   , 
negInst   ,  
SHRInst   ,  
SHRAInst  ,
SHLInst   , 
SHCInst   ,  
BrInst    ,   
BrlInst   , 
ldInst    ,  
ldrInst   ,  
stInst    ,   
strInst   ,
laInst    , 
larInst   ,
stopInst  ,
Add 		 ,
Sub 		 ,
andOp 	 ,
OrOP 		 ,
SHR 		 ,
SHRA 		 ,
SHL 		 , 
SHC 		 ,
NOTOP 	 ,
NEG 		 ,
CB 		 ,
INC4 		 ,
CONin 	 ,
Rin 		 ,
Rout 		 ,
BAout 	 ,
Gra 		 ,
Grb 		 ,
Grc 		 ,
Dec 		 ,
load 		 ,
c1out 	 ,
C2out		 ,
PCin 		 ,
PCout 	 ,
Ain 		 ,
IRin 		 ,
MDin 		 ,
MDout 	 ,
MAin 		 ,
Cout 		 ,
end_inst  ,
cpu_wait	 ,
Cin 		 ,
read_m 	 ,
write_m 	 ,
goto6 	 ,
stop		 
);

end control_unit_arch;
